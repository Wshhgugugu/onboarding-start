/*
 * Copyright (c) 2024 Shiheng
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module UWASIC_Shiheng (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  wire [7:0] en_reg_out_7_0;
  wire [7:0] en_reg_out_15_8;
  wire [7:0] en_reg_pwm_7_0;
  wire [7:0] en_reg_pwm_15_8;
  wire [7:0] pwm_duty_cycle;

  assign uio_oe = en_reg_out_15_8;

  spi_peripheral spi_peripheral_inst (
        .clk(clk),
        .rst_n(rst_n),
        .nCS(ui_in[2]),
        .SCLK(ui_in[0]),
        .COPI(ui_in[1]),
        .en_reg_out_7_0(en_reg_out_7_0),
        .en_reg_out_15_8(en_reg_out_15_8),
        .en_reg_pwm_7_0(en_reg_pwm_7_0),
        .en_reg_pwm_15_8(en_reg_pwm_15_8),
        .pwm_duty_cycle(pwm_duty_cycle)
    );

     pwm_peripheral pwm_peripheral_inst (
        .clk(clk),
        .rst_n(rst_n),
        .en_reg_out({en_reg_out_15_8, en_reg_out_7_0}),
        .en_reg_pwm({en_reg_pwm_15_8, en_reg_pwm_7_0}),
        .pwm_duty_cycle(pwm_duty_cycle),
        .pwm_out({uio_out, uo_out})
    );
    
    wire _unused = &{ui_in[7:3], uio_in, ena};

endmodule
